//for synthesis on EDA Playground
`include "DUT.sv"
`include "ALU.sv"
`include "data_mem.sv"
`include "extender.sv"
`include "instr_mem.sv"
`include "FA_1.sv"
`include "FA_4.sv"
`include "FA_8.sv"
`include "LUT_4.sv"