//effectively a 12-bit register
module PC(
         //TBD
    );

endmodule