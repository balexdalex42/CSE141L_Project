module ALU(
        input logic [7:0]   in_1, in_2,
        input 
        output logic    out_val
    );


    always_comb begin
    end
endmodule